module UART (clk, TX_D, RX_D, RTS, CTS, BYTEOUT, load);
input clk,TX_D,RTS;
output RX_D,CTS,load;
output wire [7:0]BYTEOUT;



endmodule